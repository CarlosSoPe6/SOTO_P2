module EX_MEM_PipelineRegister(
    input clk,
    input reset,
    input in_Zero,
    input in_ALUResult,
    input in_ReadData2,

    output out_Zero,
    output out_ALUResult,
    output out_ReadData2
);

endmodule // EX_MEM_PipelineRegister